//////////////////////////////////////////////////////////////////////////////////
// Company:         TSN@NNS
// Engineer:        Wenxue Wu
// 
// Create Date:     2024/05/15
// Design Name:     DFQ CAM Dequeue Process
// Module Name:     dequeue_process
// Project Name:    DFQ_CAM_v5
// Target Devices:  ZYNQ
// Tool Versions:   VIVADO 2023.2
// Description:     Dequeue process module for DFQ CAM system with FSM control
//                  Handles reading from pointer RAM and managing queue operations
// 
// Dependencies:    None
// 
// Revision:     v1.0
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module dequeue_process#(
    parameter       DATA_WIDTH = 20,
    parameter       ADDR_WIDTH = 10
)(
    input  wire                         clk,
    input  wire                         reset,
    input  wire                         start_dequeue,      // ���������ź�
    input  wire [DATA_WIDTH-1:0]        head_ptr_in,        // ��ǰ֡��ͷָ��
    input  wire [DATA_WIDTH-1:0]        ptr_ram_dout,       // ��RAM����������
    input  wire                         pcp_queue_full,     // Ŀ�����ȼ������Ƿ�����
    output reg  [ADDR_WIDTH-1:0]        ptr_ram_addr,       // �����RAM�Ķ�ȡ��ַ
    output reg  [DATA_WIDTH-1:0]        pcp_queue_din,      // ��������ȼ����е�����
    output reg                          pcp_queue_wr,       // ���ȼ����е�дʹ��
    output reg  [DATA_WIDTH-1:0]        new_head,           // ֡���Ӻ��µ�ͷָ��
    output reg                          dequeue_done,       // ֡������ɱ�־
    output reg  [15:0]                  rd_depth_cell
);

/***************function**************/

/***************parameter*************/
    localparam [3:0] ST_IDLE         = 4'd0;   // ����״̬
    localparam [3:0] ST_START        = 4'd1;   // ��ʼ����
    localparam [3:0] ST_CHECK        = 4'd2;   // ����Ƿ�Ϊβ����Ŀ
    localparam [3:0] ST_READ         = 4'd3;   // ��ȡ��������β��·����
    localparam [3:0] ST_PUSH         = 4'd4;   // �������ݵ�����
    localparam [3:0] ST_PUSH_LOOP    = 4'd5;   // ����ѭ���ȴ�
    localparam [3:0] ST_PUSH_DONE    = 4'd6;   // �������
    localparam [3:0] ST_REFRESH      = 4'd7;   // ˢ�²���
    localparam [3:0] ST_REFRESH_DONE = 4'd8;   // ˢ����ɣ�����Ƿ�Ϊָ��β��
    localparam [3:0] ST_EXIT         = 4'd9;   // �ӷ�β��·���˳�
    localparam [3:0] ST_CAM_REFRESH  = 4'd10;  // CAMˢ�²���
    localparam [3:0] ST_CAM_WAIT     = 4'd11;  // CAM�ȴ�״̬
    localparam [3:0] ST_FINAL        = 4'd12;  // ���ؿ���ǰ������״̬
    localparam [3:0] ST_EXIT2        = 4'd13;  // ��β��·���˳�
    localparam [3:0] ST_NEXT         = 4'd14;  // ��һ��������β��·����
    localparam [3:0] ST_WAIT         = 4'd15;  // �ȴ�״̬��β��·����

/***************port******************/             

/***************mechine***************/

/***************reg*******************/
    reg [3:0] current_state;
    reg [DATA_WIDTH-1:0] rd_head_reg;

/***************wire******************/
    // Flag to check if current entry is 64B (both bit 15 and 14 are set)
    wire is_cell_1 = head_ptr_in[15] && head_ptr_in[14];
    // Flag to check if current pointer entry is tail (bit 15 is set)
    wire is_last_cell = ptr_ram_dout[15];

/***************component*************/

/***************assign****************/

/***************always****************/
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            current_state    <= ST_IDLE;
            pcp_queue_wr     <= 1'b0;
            ptr_ram_addr     <= {ADDR_WIDTH{1'b0}};
            pcp_queue_din    <= {DATA_WIDTH{1'b0}};
            dequeue_done     <= 1'b0;
            new_head         <= {DATA_WIDTH{1'b0}};
            rd_head_reg      <= {DATA_WIDTH{1'b0}};
            rd_depth_cell    <= {16{1'b0}};
        end else begin
            // Default values - these signals are pulsed for one clock cycle
            pcp_queue_wr     <= 1'b0;
            dequeue_done     <= 1'b0;
            case (current_state)
                //-------------------------------------------------------------
                // State 0: IDLE - �ȴ���ʼ�ź�
                //-------------------------------------------------------------
                ST_IDLE: begin
                    if (start_dequeue) begin
                        current_state <= ST_START;
                        rd_depth_cell <= 16'b0; // Reset depth cell counter
                    end
                end

                //-------------------------------------------------------------
                // State 1: START - ��ʼ��������ͷָ��
                //-------------------------------------------------------------
                ST_START: begin
                    pcp_queue_din <= head_ptr_in;
                    pcp_queue_wr  <= 1'b1;
                    ptr_ram_addr  <= head_ptr_in[ADDR_WIDTH-1:0];
                    current_state <= ST_CHECK;
                    rd_depth_cell <= rd_depth_cell+1;
                end

                //-------------------------------------------------------------
                // State 2: CHECK - ����Ƿ�Ϊβ����Ŀ
                //-------------------------------------------------------------
                ST_CHECK: begin
                    if (is_cell_1) begin
                        current_state <= ST_EXIT;  // ��ת��β��·��
                    end else begin
                        current_state <= ST_READ;   // ������β��·��
                    end
                end

                //-------------------------------------------------------------
                // State 3: READ - ��ȡ��������β��·����
                //-------------------------------------------------------------
                ST_READ: begin
                    current_state <= ST_PUSH;
                end

                //-------------------------------------------------------------
                // State 4: PUSH - �������ݵ�����
                //-------------------------------------------------------------
                ST_PUSH: begin
                    pcp_queue_din <= ptr_ram_dout;
                    pcp_queue_wr  <= 1'b1;
                    ptr_ram_addr  <= ptr_ram_dout[ADDR_WIDTH-1:0];
                    current_state <= ST_PUSH_LOOP;
                    rd_depth_cell <= rd_depth_cell+1;
                end

                //-------------------------------------------------------------
                // State 5: PUSH_LOOP - ����ѭ���ȴ�
                //-------------------------------------------------------------
                ST_PUSH_LOOP: begin
                    current_state <= ST_PUSH_DONE;
                end

                //-------------------------------------------------------------
                // State 6: PUSH_DONE - �������
                //-------------------------------------------------------------
                ST_PUSH_DONE: begin
                    current_state <= ST_REFRESH;
                    if (is_last_cell) begin
                        ptr_ram_addr  <= ptr_ram_dout[ADDR_WIDTH-1:0];
                        current_state <= ST_EXIT;
                    end
                end

                //-------------------------------------------------------------
                // State 7: REFRESH - ˢ�²���
                //-------------------------------------------------------------
                ST_REFRESH: begin
                    current_state <= ST_REFRESH_DONE;
                    pcp_queue_din <= ptr_ram_dout;
                    ptr_ram_addr  <= ptr_ram_dout[ADDR_WIDTH-1:0];
                    pcp_queue_wr  <= 1'b1;
                    rd_depth_cell <= rd_depth_cell+1;
                end

                //-------------------------------------------------------------
                // State 8: REFRESH_DONE - ˢ����ɣ�����Ƿ�Ϊָ��β��
                //-------------------------------------------------------------
                ST_REFRESH_DONE: begin
                    if (is_last_cell) begin
                        // pcp_queue_din <= ptr_ram_dout;
                        // ptr_ram_addr  <= ptr_ram_dout[ADDR_WIDTH-1:0];
                        // pcp_queue_wr  <= 1'b1;
                        current_state <= ST_EXIT;
                    end else begin
                        current_state <= 4'd15;
                    end
                end

                4'd15: begin
                    current_state <= ST_PUSH;
                end

                //-------------------------------------------------------------
                // State 9: EXIT - �ӷ�β��·���˳�
                //-------------------------------------------------------------
                ST_EXIT: begin
                    dequeue_done  <= 1'b1;
                    current_state <= ST_CAM_REFRESH;
                end

                //-------------------------------------------------------------
                //-------------------------------------------------------------
                ST_CAM_REFRESH: begin
                    current_state <= ST_CAM_WAIT;
                    new_head      <= ptr_ram_dout;
                end

                //-------------------------------------------------------------
                // State 11: CAM_WAIT - CAM�ȴ�״̬
                //-------------------------------------------------------------
                ST_CAM_WAIT: begin
                    current_state <= ST_FINAL;
                end

                //-------------------------------------------------------------
                // State 12: FINAL - ���ؿ���ǰ������״̬
                //-------------------------------------------------------------
                ST_FINAL: begin
                    current_state <= ST_EXIT2;
                end

                ST_EXIT2: begin
                    current_state <= ST_IDLE;
                end

                //-------------------------------------------------------------
                // Default: Ĭ��״̬ - ���õ�����״̬
                //-------------------------------------------------------------
                default: begin
                    pcp_queue_wr  <= 1'b0;
                    dequeue_done  <= 1'b0;
                    current_state <= ST_IDLE;
                end
            endcase
        end
    end

endmodule